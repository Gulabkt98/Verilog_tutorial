module gate(A,B,Y);

//declaring inputs 
input A,B;
//declaring output
output Y;

//gate level modeling
//function name (port list);
//and gate (Y,A,B);
and (Y,A,B);  


endmodule